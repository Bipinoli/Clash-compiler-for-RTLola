library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.fixed_pkg.all;
use work.array_type_pkg.all;
use work.my_math_pkg.all;

--* Output Stream in the Specification
--* output trigger_gps_sats : Bool := (gps_sats.hold().defaults(to: 0) < 6)
--* Input Dependencies:
--* Storage Requirement: 0
--* Output Dependencies:
--* Stream Lookups
--* - gps_sats of Type UInt64: 0


entity trigger_gps_sats_output_stream_entity is 
	port (
		clk, pe, eval, rst : in std_logic;
			gps_sats_0 : in unsigned(63 downto 0);
			gps_sats_data_valid_0 : in std_logic;
		data_out : out bit_array(0 downto 0);
		data_valid_out : out bit_array(0 downto 0);
		pe_done_out : out std_logic;
		eval_done_out : out std_logic
	);
end trigger_gps_sats_output_stream_entity;

architecture behavioral of trigger_gps_sats_output_stream_entity is

    signal pe_done : std_logic;
    signal eval_done : std_logic;
    signal data : bit_array(0 downto 0);
    signal data_valid : bit_array(0 downto 0);

    begin

    process (clk, rst)
        -- temporal variables
		variable temp_0: unsigned(63 downto 0) := (others => '0');
		variable temp_1: unsigned(63 downto 0) := (others => '0');
		variable temp_2: unsigned(63 downto 0) := (others => '0');
		variable temp_3: unsigned(63 downto 0) := (others => '0');
		variable temp_4: std_logic := '0';
	    variable updt : std_logic := '0';
    begin
	    if (rst='1') then
	        -- Reset Phase
		    data(data'high downto 0) <= (others => '0');
		    data_valid(data_valid'high downto 0) <= (others => '0');
		    pe_done <= '0';
		    eval_done <= '0';
	    elsif (rising_edge(clk)) then
	        -- Logic Phase
	        if (pe = '1' and pe_done = '0') then
	            -- Pseudo Evaluation
                data <= data(data'high-1 downto 0) & '0';
                data_valid <= data_valid(data_valid'high-1 downto 0) & '0';
                pe_done <= '1';
		    elsif (eval = '1' and eval_done = '0') then
				-- Evaluation
				--* temp_0 := gps_sats.hold() 
				temp_0 := gps_sats_0;
				temp_1 := to_unsigned(0, 64);
				--* temp_2 := gps_sats.hold().defaults(to: 0) 
				temp_2 := sel(temp_0, temp_1, gps_sats_data_valid_0);
				temp_3 := to_unsigned(6, 64);
				--* temp_4 := (gps_sats.hold().defaults(to: 0) < 6) 
				temp_4 := to_std_logic(temp_2 < temp_3);
				updt := temp_4;
			    -- Register Update
			    data(0) <= updt;
			    data_valid(0) <= '1';
			    eval_done <= '1';
			elsif (pe = '0' and eval = '0') then
                -- Reset done Signals
                pe_done <= '0';
                eval_done <= '0';
		    end if;
	    end if;
    end process;

     -- Mapping: Register to Output Wires
    data_out <= data;
    data_valid_out <= data_valid;
    pe_done_out <= pe_done;
    eval_done_out <= eval_done;

end behavioral;
