library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.fixed_pkg.all;
use work.array_type_pkg.all;

entity hlQInterface is
    port (
        clk, rst : in std_logic;
        time_for_event : in unsigned(63 downto 0);
        time_for_deadline : in unsigned(63 downto 0);
        push_event : std_logic;
        push_deadline : in std_logic;
		x_data_in : in signed(63 downto 0);
		x_en_in : in std_logic;
		y_data_in : in signed(63 downto 0);
		y_en_in : in std_logic;
		x_data_out : out signed(63 downto 0);
		x_en_out : out std_logic;
		y_data_out : out signed(63 downto 0);
		y_en_out : out std_logic;
		a_en_out : out std_logic;
		b_en_out : out std_logic;
		c_en_out : out std_logic;
		d_en_out : out std_logic;
		e_en_out : out std_logic;
		f_en_out : out std_logic;
		g_en_out : out std_logic;
        time_out : out unsigned(63 downto 0);
        push_out : out std_logic
    );
end hlQInterface;

--* Streams and their Activation Conditions:
--* Input Streams 
--* - x @ { x }
--* - y @ { y }
--* Event-based Output Streams 
--* - a @ { x }
--* - d @ { x, y }
--* Periodic Output Streams 
--* - b @ 1000Hz
--* - c @ 2000Hz
--* - e @ 1000Hz
--* - f @ 1000Hz
--* - g @ 1000Hz
--* Resulting Deadline Array
--* || c | b, e, c, f, g ||

architecture behavioral of hlQInterface is

    -- Internal Signal Declarations
    signal clock_state_machine : integer;
    signal push_to_queue : std_logic;
	signal x_data_push : signed(63 downto 0);
	signal x_en_push: std_logic;
	signal y_data_push : signed(63 downto 0);
	signal y_en_push: std_logic;
	signal a_en_push : std_logic;
	signal b_en_push : std_logic;
	signal c_en_push : std_logic;
	signal d_en_push : std_logic;
	signal e_en_push : std_logic;
	signal f_en_push : std_logic;
	signal g_en_push : std_logic;
	signal b_en_array : bit_array(1 downto 0);
	signal c_en_array : bit_array(1 downto 0);
	signal e_en_array : bit_array(1 downto 0);
	signal f_en_array : bit_array(1 downto 0);
	signal g_en_array : bit_array(1 downto 0);
    signal last_deadline_id : integer;
    signal time_to_queue : unsigned(63 downto 0);

begin

    process(clk, rst) begin
        if (rst = '1') then
            -- Reset Phase
            clock_state_machine <= 0;
            time_to_queue <= (others => '0');
            push_to_queue <= '0';
            last_deadline_id <= 0;
			x_data_push <= (others => '0');
			x_en_push <= '0';
			y_data_push <= (others => '0');
			y_en_push <= '0';
			a_en_push <= '0';
			b_en_push <= '0';
			c_en_push <= '0';
			d_en_push <= '0';
			e_en_push <= '0';
			f_en_push <= '0';
			g_en_push <= '0';
            -- Initialize Deadline Arrays
            --* Deadline Array
            --* || c | b, e, c, f, g ||
			b_en_array(0) <= '0';
			c_en_array(0) <= '1';
			e_en_array(0) <= '0';
			f_en_array(0) <= '0';
			g_en_array(0) <= '0';
			b_en_array(1) <= '1';
			c_en_array(1) <= '1';
			e_en_array(1) <= '1';
			f_en_array(1) <= '1';
			g_en_array(1) <= '1';
        elsif (rising_edge(clk)) then
            clock_state_machine <= (clock_state_machine + 1) mod 4;
            if push_deadline = '1' and clock_state_machine = 0 then
                -- Deadline Handling
                push_to_queue <= '1';
                last_deadline_id <= (last_deadline_id + 1) mod 2;
                time_to_queue <= time_for_deadline;
				--* x @ { x }
				x_en_push <= '0';
				--* y @ { y }
				y_en_push <= '0';
				--* a @ { x }
				a_en_push <= '0';
				--* d @ { x, y }
				d_en_push <= '0';
				--* b @ 1000Hz
				b_en_push <= b_en_array(last_deadline_id);
				--* c @ 2000Hz
				c_en_push <= c_en_array(last_deadline_id);
				--* e @ 1000Hz
				e_en_push <= e_en_array(last_deadline_id);
				--* f @ 1000Hz
				f_en_push <= f_en_array(last_deadline_id);
				--* g @ 1000Hz
				g_en_push <= g_en_array(last_deadline_id);
            elsif push_event = '1' and clock_state_machine = 2 then
                -- Event Handling
                push_to_queue <= '1';
                time_to_queue <= time_for_event;
				--* x @ { x }
				x_data_push <= x_data_in;
				x_en_push <= x_en_in;
				--* y @ { y }
				y_data_push <= y_data_in;
				y_en_push <= y_en_in;
				--* a @ { x }
				a_en_push <= '1' and x_en_in;
				--* d @ { x, y }
				d_en_push <= '1' and x_en_in and y_en_in;
				--* b @ 1000Hz
				b_en_push <= '0';
				--* c @ 2000Hz
				c_en_push <= '0';
				--* e @ 1000Hz
				e_en_push <= '0';
				--* f @ 1000Hz
				f_en_push <= '0';
				--* g @ 1000Hz
				g_en_push <= '0';
            else
                -- Enable No Stream
                push_to_queue <= '0';
				x_en_push <= '0';
				y_en_push <= '0';
				a_en_push <= '0';
				b_en_push <= '0';
				c_en_push <= '0';
				d_en_push <= '0';
				e_en_push <= '0';
				f_en_push <= '0';
				g_en_push <= '0';
            end if;
        end if;
    end process;

    push_out <= push_to_queue;
    time_out <= time_to_queue;
	x_data_out <= x_data_push;
	x_en_out <= x_en_push;
	y_data_out <= y_data_push;
	y_en_out <= y_en_push;
	a_en_out <= a_en_push;
	b_en_out <= b_en_push;
	c_en_out <= c_en_push;
	d_en_out <= d_en_push;
	e_en_out <= e_en_push;
	f_en_out <= f_en_push;
	g_en_out <= g_en_push;

end behavioral;
