library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.fixed_pkg.all;
use work.array_type_pkg.all;
use work.my_math_pkg.all;

--* Output Stream in the Specification
--* output c : Int64 := (b.hold().defaults(to: 0) + b.aggregate(over: 0.1s, using: sum))
--* Input Dependencies:
--* Stream Lookups:
--* - b: 0
--* - d: 0
--* Window Lookups:
--* - d: (0.05, count)
--* Storage Requirement: 0
--* Output Dependencies:
--* Stream Lookups
--* - b of Type Int64: 0, window SlidingWin(0)
--* Window Lookups:
--* - b.aggregate(over: 0.1 s, using: sum) of type Int64


entity c_output_stream_entity is 
	port (
		clk, pe, eval, rst : in std_logic;
			b_0 : in signed(63 downto 0);
			b_data_valid_0 : in std_logic;
			b_sum_0_sw : in signed(63 downto 0);
			b_sum_0_sw_data_valid : in std_logic;
		data_out : out signed64_array(0 downto 0);
		data_valid_out : out bit_array(0 downto 0);
		pe_done_out : out std_logic;
		eval_done_out : out std_logic
	);
end c_output_stream_entity;

architecture behavioral of c_output_stream_entity is

    signal pe_done : std_logic;
    signal eval_done : std_logic;
    signal data : signed64_array(0 downto 0);
    signal data_valid : bit_array(0 downto 0);

    begin

    process (clk, rst)
        -- temporal variables
		variable temp_0: signed(63 downto 0) := (others => '0');
		variable temp_1: signed(63 downto 0) := (others => '0');
		variable temp_2: signed(63 downto 0) := (others => '0');
		variable temp_3: signed(63 downto 0) := (others => '0');
		variable temp_4: signed(63 downto 0) := (others => '0');
	    variable updt : signed(63 downto 0) := (others => '0');
    begin
	    if (rst='1') then
	        -- Reset Phase
		    data(data'high downto 0) <= (others => (others => '0'));
		    data_valid(data_valid'high downto 0) <= (others => '0');
		    pe_done <= '0';
		    eval_done <= '0';
	    elsif (rising_edge(clk)) then
	        -- Logic Phase
	        if (pe = '1' and pe_done = '0') then
	            -- Pseudo Evaluation
                data <= data(data'high-1 downto 0) & to_signed(0, updt'length);
                data_valid <= data_valid(data_valid'high-1 downto 0) & '0';
                pe_done <= '1';
		    elsif (eval = '1' and eval_done = '0') then
				-- Evaluation
				--* temp_0 := b.hold() 
				temp_0 := b_0;
				temp_1 := to_signed(0, 64);
				--* temp_2 := b.hold().defaults(to: 0) 
				temp_2 := sel(temp_0, temp_1, b_data_valid_0);
				--* temp_3 := b.aggregate(over: 0.1s, using: sum) 
				temp_3 := b_sum_0_sw;
				--* temp_4 := (b.hold().defaults(to: 0) + b.aggregate(over: 0.1s, using: sum)) 
				temp_4 := temp_2 + temp_3;
				updt := temp_4;
			    -- Register Update
			    data(0) <= updt;
			    data_valid(0) <= '1';
			    eval_done <= '1';
			elsif (pe = '0' and eval = '0') then
                -- Reset done Signals
                pe_done <= '0';
                eval_done <= '0';
		    end if;
	    end if;
    end process;

     -- Mapping: Register to Output Wires
    data_out <= data;
    data_valid_out <= data_valid;
    pe_done_out <= pe_done;
    eval_done_out <= eval_done;

end behavioral;
