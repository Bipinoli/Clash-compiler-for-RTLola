library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.fixed_pkg.all;
use work.array_type_pkg.all;
use work.my_math_pkg.all;

--* Output Stream in the Specification
--* output acceleration_x_direction_change : Bool := ((acceleration_x_rising and acceleration_x_sinking.offset(by: neg1).defaults(to: '0')) or (acceleration_x_sinking and acceleration_x_rising.offset(by: neg1).defaults(to: '0')))
--* Input Dependencies:
--* Stream Lookups:
--* - acceleration_x_changes: 
--* Window Lookups:
--* - acceleration_x_changes: (0.05, count)
--* Storage Requirement: 0
--* Output Dependencies:
--* Stream Lookups
--* - acceleration_x_rising of Type Bool: 0, -1
--* - acceleration_x_sinking of Type Bool: -1, 0


entity acceleration_x_direction_change_output_stream_entity is 
	port (
		clk, pe, eval, rst : in std_logic;
			acceleration_x_rising_0 : in std_logic;
			acceleration_x_rising_data_valid_0 : in std_logic;
			acceleration_x_rising_neg1 : in std_logic;
			acceleration_x_rising_data_valid_neg1 : in std_logic;
			acceleration_x_sinking_neg1 : in std_logic;
			acceleration_x_sinking_data_valid_neg1 : in std_logic;
			acceleration_x_sinking_0 : in std_logic;
			acceleration_x_sinking_data_valid_0 : in std_logic;
		data_out : out bit_array(0 downto 0);
		data_valid_out : out bit_array(0 downto 0);
		pe_done_out : out std_logic;
		eval_done_out : out std_logic
	);
end acceleration_x_direction_change_output_stream_entity;

architecture behavioral of acceleration_x_direction_change_output_stream_entity is

    signal pe_done : std_logic;
    signal eval_done : std_logic;
    signal data : bit_array(0 downto 0);
    signal data_valid : bit_array(0 downto 0);

    begin

    process (clk, rst)
        -- temporal variables
		variable temp_0: std_logic := '0';
		variable temp_1: std_logic := '0';
		variable temp_2: std_logic := '0';
		variable temp_3: std_logic := '0';
		variable temp_4: std_logic := '0';
		variable temp_5: std_logic := '0';
		variable temp_6: std_logic := '0';
		variable temp_7: std_logic := '0';
		variable temp_8: std_logic := '0';
		variable temp_9: std_logic := '0';
		variable temp_10: std_logic := '0';
	    variable updt : std_logic := '0';
    begin
	    if (rst='1') then
	        -- Reset Phase
		    data(data'high downto 0) <= (others => '0');
		    data_valid(data_valid'high downto 0) <= (others => '0');
		    pe_done <= '0';
		    eval_done <= '0';
	    elsif (rising_edge(clk)) then
	        -- Logic Phase
	        if (pe = '1' and pe_done = '0') then
	            -- Pseudo Evaluation
                data <= data(data'high-1 downto 0) & '0';
                data_valid <= data_valid(data_valid'high-1 downto 0) & '0';
                pe_done <= '1';
		    elsif (eval = '1' and eval_done = '0') then
				-- Evaluation
				--* temp_0 := acceleration_x_rising 
				temp_0 := acceleration_x_rising_0;
				--* temp_1 := acceleration_x_sinking.offset(by: neg1)
				temp_1 := acceleration_x_sinking_neg1;
				temp_2 := '0';
				--* temp_3 := acceleration_x_sinking.offset(by: neg1).defaults(to: '0') 
				temp_3 := sel(temp_1, temp_2, acceleration_x_sinking_data_valid_neg1);
				--* temp_4 := (acceleration_x_rising and acceleration_x_sinking.offset(by: neg1).defaults(to: '0')) 
				temp_4 := temp_0 and temp_3;
				--* temp_5 := acceleration_x_sinking 
				temp_5 := acceleration_x_sinking_0;
				--* temp_6 := acceleration_x_rising.offset(by: neg1)
				temp_6 := acceleration_x_rising_neg1;
				temp_7 := '0';
				--* temp_8 := acceleration_x_rising.offset(by: neg1).defaults(to: '0') 
				temp_8 := sel(temp_6, temp_7, acceleration_x_rising_data_valid_neg1);
				--* temp_9 := (acceleration_x_sinking and acceleration_x_rising.offset(by: neg1).defaults(to: '0')) 
				temp_9 := temp_5 and temp_8;
				--* temp_10 := ((acceleration_x_rising and acceleration_x_sinking.offset(by: neg1).defaults(to: '0')) or (acceleration_x_sinking and acceleration_x_rising.offset(by: neg1).defaults(to: '0'))) 
				temp_10 := temp_4 or temp_9;
				updt := temp_10;
			    -- Register Update
			    data(0) <= updt;
			    data_valid(0) <= '1';
			    eval_done <= '1';
			elsif (pe = '0' and eval = '0') then
                -- Reset done Signals
                pe_done <= '0';
                eval_done <= '0';
		    end if;
	    end if;
    end process;

     -- Mapping: Register to Output Wires
    data_out <= data;
    data_valid_out <= data_valid;
    pe_done_out <= pe_done;
    eval_done_out <= eval_done;

end behavioral;
